/*
 * Stack_test.cpp
 *
 *  Created on: Feb 13, 2021
 *      Author: abdulwaheed
 */

#include "Stack.h"

int main() {
	return 0;
}
